.title KiCad schematic
.include "models/BZX84C4V7.spice.txt"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/C2012CH2A103J125AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C3225X7S1H106M250AB_p.mod"
.include "models/US1M.spice.txt"
.include "models/ZXCT1030.spice.txt"
.include "models/ZXMN3B14F.spice.txt"
.include "models/ZXMP3A17E6.spice.txt"
V1 /VIN 0 20
V2 +5V 0 5
XU2 +5V 0 C3225X7S1H106M250AB_p
XU3 +5V 0 C2012X7R2A104K125AA_p
R1 /VIN /OCP 0.47
XU4 /VIN /VSN C2012C0G2A102J060AA_p
R4 /OCP /VSN 10k
R5 +5V /COMP_OUT 68k
R3 /OCP /DRAIN 4.7K
R7 /CURRENT_FEEDBACK /VOCM 120
XU8 /CURRENT_FEEDBACK 0 C2012CH2A103J125AA_p
XU7 0 /CURRENT_FEEDBACK DI_BZX84C4V7
XU6 +5V /VSN /VIN 0 /TRP NC_01 /VOCM /COMP_OUT ZXCT1030
R9 +5V /TRP 9.76k
R11 /TRP 0 8.66k
XU1 /VOUT /DRAIN /OCP ZXMP3A17E6
XU5 /DRAIN /GATE 0 ZXMN3B14F
R12 /VOUT 0 50
R2 /VIN /OCP 0.47
R6 /COMP_OUT /GATE 10
D1 /GATE /COMP_OUT DI_US1M
.end
